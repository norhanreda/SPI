module Master(clk, reset,start, slaveSelect, masterDataToSend, masterDataReceived,SCLK, CS, MOSI, MISO);
input  wire clk; // Clock which is sent from the testbench to the master.
input wire reset; // Reset which is sent from the testbench to all the modules.
input wire start; // This signals the master to start the transmission (also the master will read "masterDataToSend" in order to send it to the slave).
input wire [1:0] slaveSelect; // This tells the master which slave to transmit to. It should be read by the master when "start" becomes high.
input wire [7:0] masterDataToSend; // What data should the master send to the slave during the transmission
output reg [7:0] masterDataReceived; // What data did the master receive from the slave during the past transmission
output reg SCLK; // The clock generated by the master for the transmission. The master uses the "clk" to generate this signal. Both the master and the slave can only use this signal for synchronizing the transmission. 
output reg  [0:2] CS; // The chip select signal used by the master to select a slave. If a slave is selected, the master should set its corresponding CS to 0 (active low).
output reg MOSI; // The data signal going from the master to the slave.
input wire  MISO; // The data signal going from the slave to the master.

reg [7:0] t_reg;
integer count;
always @(slaveSelect)
begin
case (slaveSelect)
       2'b00:CS=3'b011;
       2'b 01: CS=3'b101;   
       2'b10: CS=3'b110;
 
      default: CS=3'b111;
    endcase
end 
always @(posedge reset)
begin 
count<=-1;
t_reg<=8'b00000000;
 MOSI<=0;
masterDataReceived<=8'b00000000;
end
always #5 SCLK=~clk;
always @( posedge start )//
begin
t_reg<=masterDataToSend;
count<=0;
end
always @(posedge  SCLK)//sending
begin 
if(reset==0)begin
if((CS[0]==0) || (CS[1]==0) || (CS[2]==0) )
begin
if(count>=0 && count<=8)//7-8

begin
MOSI<=t_reg[7];
end

if(count==9) 
begin
count<=-1;
end
end
if((CS[0]==1) && (CS[1]==1) && (CS[2]==1) )
MOSI<=1'bz;
end
end 
///////////////////////////////////////////
always @ (negedge SCLK)
begin
if(reset==0)begin
if((CS[0]==0) || (CS[1]==0) || (CS[2]==0) )
 
begin
if(count>=0 && count<=8)
begin

t_reg<=t_reg<<<1;
t_reg[0]<=0;
t_reg[0]<=MISO;
count=count+1;
end
end
if(count==9)
begin
masterDataReceived<=t_reg;
count<=-1;

end
end
end 
endmodule
